module top (

);

endmodule


module uart_sim (
    input clk,
    input rst,
    input rx_i,
    output tx_o
);

top #() top_uut (.*);

endmodule
